signal d0_0: std_logic_vector(15 downto 0);
signal d0_1: std_logic_vector(15 downto 0);
signal d0_2: std_logic_vector(14 downto 0);
signal d0_3: std_logic_vector(12 downto 0);
signal d0_4: std_logic_vector(11 downto 0);
signal d1_0: std_logic_vector(15 downto 0);
signal d1_1: std_logic_vector(15 downto 0);
signal d1_2: std_logic_vector(14 downto 0);
signal d1_3: std_logic_vector(13 downto 0);
signal d2_0: std_logic_vector(15 downto 0);
signal d2_1: std_logic_vector(15 downto 0);
signal d2_2: std_logic_vector(15 downto 0);
