signal d0_0: std_logic_vector(47 downto 0);
signal d0_1: std_logic_vector(47 downto 0);
signal d0_2: std_logic_vector(46 downto 0);
signal d0_3: std_logic_vector(44 downto 0);
signal d0_4: std_logic_vector(42 downto 0);
signal d0_5: std_logic_vector(40 downto 0);
signal d0_6: std_logic_vector(38 downto 0);
signal d0_7: std_logic_vector(36 downto 0);
signal d0_8: std_logic_vector(34 downto 0);
signal d0_9: std_logic_vector(32 downto 0);
signal d0_10: std_logic_vector(30 downto 0);
signal d0_11: std_logic_vector(28 downto 0);
signal d0_12: std_logic_vector(27 downto 0);
signal d1_0: std_logic_vector(47 downto 0);
signal d1_1: std_logic_vector(47 downto 0);
signal d1_2: std_logic_vector(46 downto 0);
signal d1_3: std_logic_vector(44 downto 0);
signal d1_4: std_logic_vector(42 downto 0);
signal d1_5: std_logic_vector(40 downto 0);
signal d1_6: std_logic_vector(38 downto 0);
signal d1_7: std_logic_vector(36 downto 0);
signal d1_8: std_logic_vector(35 downto 0);
signal d2_0: std_logic_vector(47 downto 0);
signal d2_1: std_logic_vector(47 downto 0);
signal d2_2: std_logic_vector(46 downto 0);
signal d2_3: std_logic_vector(44 downto 0);
signal d2_4: std_logic_vector(42 downto 0);
signal d2_5: std_logic_vector(41 downto 0);
signal d3_0: std_logic_vector(47 downto 0);
signal d3_1: std_logic_vector(47 downto 0);
signal d3_2: std_logic_vector(46 downto 0);
signal d3_3: std_logic_vector(45 downto 0);
signal d4_0: std_logic_vector(47 downto 0);
signal d4_1: std_logic_vector(47 downto 0);
signal d4_2: std_logic_vector(47 downto 0);
